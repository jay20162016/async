`include "delay_one.sv"
`include "delay.sv"
`include "delay_multi.sv"

`include "hlatch.sv"

`include "source.sv"
`include "sink.sv"

`include "split.sv"
`include "combine.sv"

`include "merge.sv"
`include "merge2.sv"

`include "mux.sv"
`include "mux2.sv"

`include "demux.sv"
`include "demux2.sv"

`include "cond_sink.sv"
`include "cond_sink2.sv"

`include "mutex.sv"
`include "arbiter.sv"
