(* blackbox, keep *)
module loop_breaker(input A, output Y);
  assign Y = A;
endmodule
