// does not include common/*
`include "delay/delay_one.sv"
`include "delay/delay.sv"
`include "delay/delay_multi.sv"

`include "active/hlatch.sv"

`include "active/source.sv"
`include "active/sink.sv"

`include "flow/split.sv"
`include "flow/combine.sv"

`include "flow/merge.sv"
`include "flow/merge2.sv"

`include "condflow/mux.sv"
`include "condflow/mux2.sv"

`include "condflow/demux.sv"
`include "condflow/demux2.sv"

`include "condflow/cond_sink.sv"
`include "condflow/cond_sink2.sv"

`include "condflow/swap.sv"
`include "condflow/swap2.sv"

`include "condflow/swap_sink.sv"
`include "condflow/swap_sink2.sv"

`include "arbiter/mutex.sv"
`include "arbiter/arbiter.sv"

`include "logic/and.sv"
`include "logic/xor.sv"

`include "arith/add1.sv"
