`include "delay_one.v"
`include "delay.v"
`include "delay_multi.v"

`include "hlatch.v"

`include "source.v"
`include "sink.v"

`include "split.v"
`include "combine.v"

`include "merge.v"
`include "merge2.v"

`include "mux.v"
`include "mux2.v"

`include "demux.v"
`include "demux2.v"

`include "cond_sink.v"
`include "cond_sink2.v"

`include "mutex.v"
`include "arbiter.v"
